`include "ram_mod.v"
`include "cache_mod.v"

module cache_and_ram #(parameter cache_index_size=5)(
	
);








ram_mod ram();
cache_mod cache();
	

	

endmodule 
